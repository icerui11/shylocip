    �   <��I �d�      �        �I  �I$�I$I$� �I$��I  �$�I$�@ � �?�I$�@ � > � � � � �UPP�� z � � � � � � � � �� �s��!BP�BB����� �!!BB�!�""!" ��D@ � 7�� �@�DD�D!���B�D � � �    �@ �" �!A" � � ���� {����� �B" � �B � � � � � � �B! �~�ǄB�! �!B  > �B� ��BABA0�D  |�? �  �A �!��}���a� �A!�  � ��A z�  �$!AA�}�$!ABA��BA" � > ���� �HB� � � ���?��!A ��q�� � � > � > � ?�?� �A�>�8!��$AA �AAA @� ��?�� ~@��@�! A��}�pA ���P� �! @�@��� � � ���P� A =������ ������ �A @؄ � �  � � v ހ� ;� �>���� �A D  � 7�� ���?�>��AA @�	!� 8��y$D � A� @�"! �� � �   6� ��`� ��  �B A  �        