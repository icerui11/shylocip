             