        <��I �d�  �� ����/����`  �� M���6�wĜ��� _� �x� nz?�����` ��
v�G!ܥ s�� � �bF 1�i��2   -�  q�  �Vx�1�y��� ��1F]?/�[?���  >��  ��
P���}� h +cn9���   S�����/6E�}� k�� ���O ��r�� ��4  BȀ ��"U��� $�  H�� ��"�4�
߀ _`�܇h�5�� ����̰����� � �P 4� ]�U���  G� � �-3��cJ����_H��?��b��F����w m�@ Z�>(�]�(�+㎀C7`?�pXB���qD��0��=�Ie����^�&ڢ9]�i'b���>)�����2LX�D"��c$��6����r?7a��On�9��=�5o[����pN�}��8E-s�?����-ip@�p;���!`�8�?-�(Nz(AK�^z�x}AFN}H�ҐJJG=A�g�|��^ ��n���bD0]�C�S��̬�4��.���<F��C���?p��B��<"��#X�/�"�����.��d��Rd�IrhD����clʎ~�aq��R�RG����s�_�!i�������'�ɕg��7ނx�*@��,)��)��4��ɺ�`���A�e%
:.#�����^tw��h͙�v�EÁ��W�����aa�X�ک�qWK�:�����_1&��K�����=�$�S)���/��;��*Ώ��7��Z$?_�8�N�E����o@��Y�5�E��Ta,�F�ak�a�4ESanPk:�DV��\�_���&�NG-��;���-(�6/&�r���|��B���C!�R�1J\�r�h?��SF
j��qy�<Ѽ��3�)a���:��(_�%�C���I��52\n�=?��;(Q).��D�V�ٳ���0q�j���Y��_�<��<id�"��O�J��QKT�zG�R�iL ���J��M�W�G���(F�<��C�Y����H]%غ>���?�w9	�"���4f2��_1u�I��V1�(\��e��8���`��?��Bu0��d��/rZ�>��H47������qH�{j3r�n�䡡@팘�Zd0߈�����:H��:������K�6Y;��~qh���Z�Q4q�;��eh�jMSϱ����*<��Ay�1�&0�:3�r���?��<��v�_D~�'�L$�|�����"'͞��)����t\��X	��ա����G�)��[���z�ǯ��� =����0�p/�	�,�&�I��ӄ�
	հP�/(f٢���x�j	�j�>�"
s���DXX2=O�z�� �#VBL��ux�)�oM�؁��!���T7K���z��.#p����7\3kȘ�T"5�FFۡ%X�/��\�q�D�����7��"/���왯 F��)3�1��sP�əν���"5j� �"�dй6:.�,�lf����nդ��xˠ�8b��´��bg6K�#� ��7������2*���u�Ѹ�񅖹�P3�V�H�/f5	sF-��f�@��������l���\�G[�k���'e2�i�HR������ڄ�A)�uj"����K�F}W0��v�m�nQ�IQe��d1��X?������p�7����Iq��ہ�yl�`R��k�����f����"?����!� q�<����� f�dĈ��x�$�EHP�$�$�XJy$���d�s8t\�E�q,(]�ߎ�ù@�*0��BA����_�Ӫ�7�,"3xO����<)#0����n!��3���Xp��K���FA関��qf��a�C�`���Ѳ?��I�v?����v�Qǁ�L?�)�#�T�b��Tr�`�2F�)�>���㑐��]^`!B�I�R��6i�[�"G9���Mc��h���&׉٣�H���-2c���|��.D��'ؒ.Z�y     